module mctrl_tb();

endmodule